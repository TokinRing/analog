module init_const (
constant);

output [7:0] constant;
reg [7:0] constant;

always	
	constant = 8'b10000000;
	
endmodule